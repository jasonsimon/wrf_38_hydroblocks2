    Mac OS X            	   2  �     �                                      ATTR      �   �  P                  �  P  #com.apple.fileutil.PlaceholderData   DENO      P                     0          �      d7eb0e052603423e9295380800f0914e        d7eb0e052603423e9295380800f0914e        1e46c45d49c44968881c65a8ad8230a3        bbcf29b55b6743d9966ac394017d2878        7a8eae03921e40b0b276dd4fcb35374a                                                aa515e15-a5b2-4b80-9555-0e9535c7e498   